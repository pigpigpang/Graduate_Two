library IEEE;
use IEEE.STD_LOGIC_1164.all;
entity decoder38 is
port( a:in STD_LOGIC_VECTOR(2 downto 0);
	  q:out STD_LOGIC_VECTOR(7 downto 0));
end decoder38 ;
architecture decoder38_arch of decoder38 is
begin
	process(a)
	begin
		case a is
			when "000" =>q<="00000001";
			when "001" =>q<="00000010";
			when "010" =>q<="00000100";
			when "011" =>q<="00001000";
			when "100" =>q<="00010000";
			when "101" =>q<="00100000";
			when "110" =>q<="01000000";
			when "111" =>q<="10000000";
			when others =>null;
		end case;
	end process;
end decoder38_arch;	